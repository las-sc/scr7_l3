
// Flits signal widths
// REQ
parameter   SCR_BASE_CL3_NOC_REQ_OPC_WIDTH      =   7;
parameter   SCR_BASE_CL3_NOC_DAT_DATAID_WIDTH   =   2;
parameter   SCR_BASE_CL3_NOC_REQ_SIZE_WIDTH     =   3;
parameter   SCR_BASE_CL3_NOC_REQ_PCTYPE_WIDTH   =   4;
parameter   SCR_BASE_CL3_NOC_REQ_MEMATTR_WIDTH  =   4;
parameter   SCR_BASE_CL3_NOC_REQ_SNPATTR_WIDTH  =   1;
parameter   SCR_BASE_CL3_NOC_REQ_EXCL_WIDTH     =   1;

// RSP
parameter   SCR_BASE_CL3_NOC_RSP_OPC_WIDTH      =   5;
parameter   SCR_BASE_CL3_NOC_RSP_RESPERR_WIDTH  =   2;
parameter   SCR_BASE_CL3_NOC_RSP_RESP_WIDTH     =   3;
parameter   SCR_BASE_CL3_NOC_RSP_PCTYPE_WIDTH   =   4;

// SNP
parameter   SCR_BASE_CL3_NOC_SNP_OPC_WIDTH      =   5;
parameter   SCR_BASE_CL3_NOC_SNP_RTOSRC_WIDTH   =   1;

// DAT
parameter   SCR_BASE_CL3_NOC_DAT_OPC_WIDTH      =   4;
parameter   SCR_BASE_CL3_NOC_DAT_RESPERR_WIDTH  =   2;
parameter   SCR_BASE_CL3_NOC_DAT_RESP_WIDTH     =   3;
parameter   SCR_BASE_CL3_NOC_DAT_FSTATE_WIDTH   =   4;
parameter   SCR_BASE_CL3_NOC_DAT_CCID_WIDTH     =   2;

// REQ Flits
parameter   [SCR_BASE_CL3_NOC_REQ_OPC_WIDTH-1:0]    SCR_BASE_CHI_REQ_READSHARED             = 'h1;
parameter   [SCR_BASE_CL3_NOC_REQ_OPC_WIDTH-1:0]    SCR_BASE_CHI_REQ_READCLEAD              = 'h2;
parameter   [SCR_BASE_CL3_NOC_REQ_OPC_WIDTH-1:0]    SCR_BASE_CHI_REQ_READONCE               = 'h3;
parameter   [SCR_BASE_CL3_NOC_REQ_OPC_WIDTH-1:0]    SCR_BASE_CHI_REQ_READNOSNP              = 'h4;
parameter   [SCR_BASE_CL3_NOC_REQ_OPC_WIDTH-1:0]    SCR_BASE_CHI_REQ_READUNIC               = 'h7;
parameter   [SCR_BASE_CL3_NOC_REQ_OPC_WIDTH-1:0]    SCR_BASE_CHI_REQ_CLEANSHARED            = 'h8;
parameter   [SCR_BASE_CL3_NOC_REQ_OPC_WIDTH-1:0]    SCR_BASE_CHI_REQ_CLEANINVALID           = 'h9;
parameter   [SCR_BASE_CL3_NOC_REQ_OPC_WIDTH-1:0]    SCR_BASE_CHI_REQ_MAKEINVALID            = 'ha;
parameter   [SCR_BASE_CL3_NOC_REQ_OPC_WIDTH-1:0]    SCR_BASE_CHI_REQ_CLEANUNIC              = 'hb;
parameter   [SCR_BASE_CL3_NOC_REQ_OPC_WIDTH-1:0]    SCR_BASE_CHI_REQ_MAKEUNIC               = 'hc;
parameter   [SCR_BASE_CL3_NOC_REQ_OPC_WIDTH-1:0]    SCR_BASE_CHI_REQ_EVICT                  = 'hd;
parameter   [SCR_BASE_CL3_NOC_REQ_OPC_WIDTH-1:0]    SCR_BASE_CHI_REQ_READNOSNPSEP           = 'h11;
parameter   [SCR_BASE_CL3_NOC_REQ_OPC_WIDTH-1:0]    SCR_BASE_CHI_REQ_WRITEEVICTFULL         = 'h15;
parameter   [SCR_BASE_CL3_NOC_REQ_OPC_WIDTH-1:0]    SCR_BASE_CHI_REQ_WRITECLEANFULL         = 'h17;
parameter   [SCR_BASE_CL3_NOC_REQ_OPC_WIDTH-1:0]    SCR_BASE_CHI_REQ_WRITEUNICPTL           = 'h18;
parameter   [SCR_BASE_CL3_NOC_REQ_OPC_WIDTH-1:0]    SCR_BASE_CHI_REQ_WRITEUNICFULL          = 'h19;
parameter   [SCR_BASE_CL3_NOC_REQ_OPC_WIDTH-1:0]    SCR_BASE_CHI_REQ_WRITEBACKPTL           = 'h1a;
parameter   [SCR_BASE_CL3_NOC_REQ_OPC_WIDTH-1:0]    SCR_BASE_CHI_REQ_WRITEBACKFULL          = 'h1b;
parameter   [SCR_BASE_CL3_NOC_REQ_OPC_WIDTH-1:0]    SCR_BASE_CHI_REQ_WRITENOSNPPTL          = 'h1c;
parameter   [SCR_BASE_CL3_NOC_REQ_OPC_WIDTH-1:0]    SCR_BASE_CHI_REQ_WRITENOSNPFULL         = 'h1d;
parameter   [SCR_BASE_CL3_NOC_REQ_OPC_WIDTH-1:0]    SCR_BASE_CHI_REQ_READONCECLEANINVALID   = 'h24;
parameter   [SCR_BASE_CL3_NOC_REQ_OPC_WIDTH-1:0]    SCR_BASE_CHI_REQ_READONCEMAKEINVALID    = 'h25;
parameter   [SCR_BASE_CL3_NOC_REQ_OPC_WIDTH-1:0]    SCR_BASE_CHI_REQ_READNOTSHAREDDIRTY     = 'h26;
parameter   [SCR_BASE_CL3_NOC_REQ_OPC_WIDTH-1:0]    SCR_BASE_CHI_REQ_CLEANSHAREDPERSIST     = 'h27;
parameter   [SCR_BASE_CL3_NOC_REQ_OPC_WIDTH-1:0]    SCR_BASE_CHI_REQ_MAKEREADUNIC           = 'h41;
parameter   [SCR_BASE_CL3_NOC_REQ_OPC_WIDTH-1:0]    SCR_BASE_CHI_REQ_WRITEEVICTOREVICT      = 'h42;
parameter   [SCR_BASE_CL3_NOC_REQ_OPC_WIDTH-1:0]    SCR_BASE_CHI_REQ_WRITEUNICZERO          = 'h43;
parameter   [SCR_BASE_CL3_NOC_REQ_OPC_WIDTH-1:0]    SCR_BASE_CHI_REQ_WRITENOSNPZERO         = 'h44;
parameter   [SCR_BASE_CL3_NOC_REQ_OPC_WIDTH-1:0]    SCR_BASE_CHI_REQ_READPREFERUNIC         = 'h4c;
parameter   [SCR_BASE_CL3_NOC_REQ_OPC_WIDTH-1:0]    SCR_BASE_CHI_REQ_WRITENOSNPFULLCLEANSH  = 'h50;
parameter   [SCR_BASE_CL3_NOC_REQ_OPC_WIDTH-1:0]    SCR_BASE_CHI_REQ_WRITENOSNPFULLCLEANINV = 'h51;
parameter   [SCR_BASE_CL3_NOC_REQ_OPC_WIDTH-1:0]    SCR_BASE_CHI_REQ_WRITENOSNPFULLCLEANSHPERSEP    = 'h52;
parameter   [SCR_BASE_CL3_NOC_REQ_OPC_WIDTH-1:0]    SCR_BASE_CHI_REQ_WRITEUNICFULLCLEANSH   = 'h54;
parameter   [SCR_BASE_CL3_NOC_REQ_OPC_WIDTH-1:0]    SCR_BASE_CHI_REQ_WRITEUNICFULLCLEANSHPERSEP     = 'h56;
parameter   [SCR_BASE_CL3_NOC_REQ_OPC_WIDTH-1:0]    SCR_BASE_CHI_REQ_WRITEBACKFULLCLEANSH   = 'h58;
parameter   [SCR_BASE_CL3_NOC_REQ_OPC_WIDTH-1:0]    SCR_BASE_CHI_REQ_WRITEBACKFULLCLEANINV  = 'h59;
parameter   [SCR_BASE_CL3_NOC_REQ_OPC_WIDTH-1:0]    SCR_BASE_CHI_REQ_WRITEBACKFULLCLEANSHPERSEP     = 'h5a;
parameter   [SCR_BASE_CL3_NOC_REQ_OPC_WIDTH-1:0]    SCR_BASE_CHI_REQ_WRITECLEANFULLCLEANSH  = 'h5c;
parameter   [SCR_BASE_CL3_NOC_REQ_OPC_WIDTH-1:0]    SCR_BASE_CHI_REQ_WRITECLEANFULLCLEANSHPERSEP    = 'h5e;
parameter   [SCR_BASE_CL3_NOC_REQ_OPC_WIDTH-1:0]    SCR_BASE_CHI_REQ_WRITENOSNPPTLCLEANSH   = 'h60;
parameter   [SCR_BASE_CL3_NOC_REQ_OPC_WIDTH-1:0]    SCR_BASE_CHI_REQ_WRITENOSNPPTLCLEANINV  = 'h61;
parameter   [SCR_BASE_CL3_NOC_REQ_OPC_WIDTH-1:0]    SCR_BASE_CHI_REQ_WRITENOSNPPTLCLEANSHPERSEP     = 'h62;
parameter   [SCR_BASE_CL3_NOC_REQ_OPC_WIDTH-1:0]    SCR_BASE_CHI_REQ_WRITEUNICPTLCLEANSH    = 'h64;
parameter   [SCR_BASE_CL3_NOC_REQ_OPC_WIDTH-1:0]    SCR_BASE_CHI_REQ_WRITEUNICPTLCLEANSHPERSEP      = 'h66;

// RSP Flits
parameter   [SCR_BASE_CL3_NOC_RSP_OPC_WIDTH-1:0]    SCR_BASE_CHI_RSP_SNPRESP                = 'h1;
parameter   [SCR_BASE_CL3_NOC_RSP_OPC_WIDTH-1:0]    SCR_BASE_CHI_RSP_COMPACK                = 'h2;
parameter   [SCR_BASE_CL3_NOC_RSP_OPC_WIDTH-1:0]    SCR_BASE_CHI_RSP_COMP                   = 'h4;
parameter   [SCR_BASE_CL3_NOC_RSP_OPC_WIDTH-1:0]    SCR_BASE_CHI_RSP_COMPDBIDRESP           = 'h5;
parameter   [SCR_BASE_CL3_NOC_RSP_OPC_WIDTH-1:0]    SCR_BASE_CHI_RSP_DBIDRESP               = 'h6;
parameter   [SCR_BASE_CL3_NOC_RSP_OPC_WIDTH-1:0]    SCR_BASE_CHI_RSP_READRECEIPT            = 'h8;
parameter   [SCR_BASE_CL3_NOC_RSP_OPC_WIDTH-1:0]    SCR_BASE_CHI_RSP_SNPRESPFWDED           = 'h9;
parameter   [SCR_BASE_CL3_NOC_RSP_OPC_WIDTH-1:0]    SCR_BASE_CHI_RSP_RESPSEPDATA            = 'hb;
parameter   [SCR_BASE_CL3_NOC_RSP_OPC_WIDTH-1:0]    SCR_BASE_CHI_RSP_PERSIST                = 'hc;
parameter   [SCR_BASE_CL3_NOC_RSP_OPC_WIDTH-1:0]    SCR_BASE_CHI_RSP_COMPPERSIST            = 'hd;
parameter   [SCR_BASE_CL3_NOC_RSP_OPC_WIDTH-1:0]    SCR_BASE_CHI_RSP_DBIDRESPORD            = 'he;

// SNP Flits
parameter   [SCR_BASE_CL3_NOC_SNP_OPC_WIDTH-1:0]    SCR_BASE_CHI_SNP_SNPSHARED              = 'h1;
parameter   [SCR_BASE_CL3_NOC_SNP_OPC_WIDTH-1:0]    SCR_BASE_CHI_SNP_SNPCLEAN               = 'h2;
parameter   [SCR_BASE_CL3_NOC_SNP_OPC_WIDTH-1:0]    SCR_BASE_CHI_SNP_SNPONCE                = 'h3;
parameter   [SCR_BASE_CL3_NOC_SNP_OPC_WIDTH-1:0]    SCR_BASE_CHI_SNP_SNPNOTSHAREDDIRTY      = 'h4;
parameter   [SCR_BASE_CL3_NOC_SNP_OPC_WIDTH-1:0]    SCR_BASE_CHI_SNP_SNPUNIC                = 'h7;
parameter   [SCR_BASE_CL3_NOC_SNP_OPC_WIDTH-1:0]    SCR_BASE_CHI_SNP_SNPCLEANSHARED         = 'h8;
parameter   [SCR_BASE_CL3_NOC_SNP_OPC_WIDTH-1:0]    SCR_BASE_CHI_SNP_SNPCLEANINVALID        = 'h9;
parameter   [SCR_BASE_CL3_NOC_SNP_OPC_WIDTH-1:0]    SCR_BASE_CHI_SNP_SNPMAKEINVALID         = 'ha;
parameter   [SCR_BASE_CL3_NOC_SNP_OPC_WIDTH-1:0]    SCR_BASE_CHI_SNP_SNPSHAREDFWD           = 'h11;
parameter   [SCR_BASE_CL3_NOC_SNP_OPC_WIDTH-1:0]    SCR_BASE_CHI_SNP_SNPCLEANFWD            = 'h12;
parameter   [SCR_BASE_CL3_NOC_SNP_OPC_WIDTH-1:0]    SCR_BASE_CHI_SNP_SNPONCEFWD             = 'h13;
parameter   [SCR_BASE_CL3_NOC_SNP_OPC_WIDTH-1:0]    SCR_BASE_CHI_SNP_SNPNOTSHAREDDIRTYFWD   = 'h14;
parameter   [SCR_BASE_CL3_NOC_SNP_OPC_WIDTH-1:0]    SCR_BASE_CHI_SNP_SNPPREFERUNIC          = 'h15;
parameter   [SCR_BASE_CL3_NOC_SNP_OPC_WIDTH-1:0]    SCR_BASE_CHI_SNP_SNPPREFERUNICFWD       = 'h16;
parameter   [SCR_BASE_CL3_NOC_SNP_OPC_WIDTH-1:0]    SCR_BASE_CHI_SNP_SNPUNICFWD             = 'h17;

// DAT Flits
parameter   [SCR_BASE_CL3_NOC_DAT_OPC_WIDTH-1:0]    SCR_BASE_CHI_DAT_OPC_SNPRESPDATA        = 'h1;
parameter   [SCR_BASE_CL3_NOC_DAT_OPC_WIDTH-1:0]    SCR_BASE_CHI_DAT_COPYBACKWRDATA         = 'h2;
parameter   [SCR_BASE_CL3_NOC_DAT_OPC_WIDTH-1:0]    SCR_BASE_CHI_DAT_NONCOPYBACKWRDATA      = 'h3;
parameter   [SCR_BASE_CL3_NOC_DAT_OPC_WIDTH-1:0]    SCR_BASE_CHI_DAT_COMPDATA               = 'h4;
parameter   [SCR_BASE_CL3_NOC_DAT_OPC_WIDTH-1:0]    SCR_BASE_CHI_DAT_SNPRESPDATAPTL         = 'h5;
parameter   [SCR_BASE_CL3_NOC_DAT_OPC_WIDTH-1:0]    SCR_BASE_CHI_DAT_SNPRESPDATAFWDED       = 'h6;
parameter   [SCR_BASE_CL3_NOC_DAT_OPC_WIDTH-1:0]    SCR_BASE_CHI_DAT_WRITEDATACANCEL        = 'h7;
parameter   [SCR_BASE_CL3_NOC_DAT_OPC_WIDTH-1:0]    SCR_BASE_CHI_DAT_DATASEPRESP            = 'hb;
parameter   [SCR_BASE_CL3_NOC_DAT_OPC_WIDTH-1:0]    SCR_BASE_CHI_DAT_NCBWRDATACOMPACK       = 'hc;


endpackage: scr_base_cl3_chipkg
