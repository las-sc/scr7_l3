///
/// @file       <scr_base_l3_bk_filelist.sv>
/// @brief      L3 Bank File List
/// @author     esk-sc
///
/// Copyright by Syntacore LLC (C) (2016 - 2021). ALL RIGHTS RESERVED. STRICTLY CONFIDENTIAL.
/// Information contained in this material is confidential and propri
/// and its affiliates and may not be modified, copied, published, di
/// displayed or exhibited, in either electronic or printed formats w
/// authorization of the Syntacore LLC. Subject to License Agreement.

// Parameters and Macros
`include "scr_base_int_description.svh"
`include "scr_base_l3_default_config.svh"

`include "scr_base_cl3_chipkg.sv"

`include "scr_base_l3_funcs_pkg.sv"
`include "scr_base_l3_params_pkg.sv"
`include "scr_base_l3_types_pkg.sv"

`include "scr_base_l3_description.svh"

// Submodules
`include "scr_base_l3_bk_dp.sv"
`include "scr_base_l3_bk_rob.sv"
`include "scr_base_l3_bk_tp.sv"
`include "scr_base_l3_bk.sv"
