`ifndef __SCR_BASE_INT_DESCRIPTION_DEFINED__
`define __SCR_BASE_INT_DESCRIPTION_DEFINED__
///
/// @file     <scr_base_int_description.svh>
/// @brief    Internal Architecture Description file
/// @authors  esk-sc
///
/// Copyright by Syntacore LLC (C) (2016 - 2021). ALL RIGHTS RESERVED. STRICTLY CONFIDENTIAL.
/// Information contained in this material is confidential and proprietary to Syntacore LLC
/// and its affiliates and may not be modified, copied, published, disclosed, distributed,
/// displayed or exhibited, in either electronic or printed formats without written
/// authorization of the Syntacore LLC. Subject to License Agreement.
///

`include "scr_base_l3_default_config.svh"

`endif // __SCR_BASE_INT_DESCRIPTION_DEFINED__
