`ifndef __SCR_BASE_L3_DESCRITION_DEFINED__
`define __SCR_BASE_L3_DESCRITION_DEFINED__
///
/// @file       <scr_base_l3_params.svh>
/// @brief      L3$ Parameters declaration
///
/// @authors    esk-sc
////
/// Copyright by Syntacore LLC (C) (2016 - 2021). ALL RIGHTS RESERVED. STRICTLY CONFIDENTIAL.
/// Information contained in this material is confidential and proprietary to Syntacore LLC
/// and its affiliates and may not be modified, copied, published, disclosed, distributed,
/// displayed or exhibited, in either electronic or printed formats without written
/// authorization of the Syntacore LLC. Subject to License Agreement.
///






`endif //__SCR_BASE_L3_DESCRITION_DEFINED__